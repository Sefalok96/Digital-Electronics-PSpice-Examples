
V1 N001 0 15v
V2 0 N004 10v
R1 N001 N002 10k
R2 N003 N004 5k
D1 N002 0 DA
D2 N002  N003 DA

.model DA D(Ron=0.0001 Roff=100G Vfwd=0)
.lib C:\Users\Sefa\Desktop\Library\lib.txt
.tran 20m
.backanno
.end
