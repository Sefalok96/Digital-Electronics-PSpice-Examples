
Vin N001 0 PULSE(0 5 0 0 0 1m 5m)
C N003 N004 1u
R N004 N005 6.8k
VD N005 0 5V
X1 N001 N002 N003 N005 0 CD4001
X2 N004 N004 N002 N005 0 CD4001

.lib C:\Users\Sefa\Desktop\Library\Digilib.txt
.tran 20m
.backanno
.end